// Multiplexer

module Mux(sel, A1, B1, Mux_out);

input sel;
input [31:0] A1, B1;
output [31:0] Mux_out;

assign Mux_out = (sel==1'b0) ? A1 : B1;

endmodule